module bcdex3(x,y);
input [3:0]x;
output [3:0]y;
assign y=x+4'b0011;
endmodule



